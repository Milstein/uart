`timescale 1ns / 1ps
module transmitter
(
	input wire [7:0] din,
	input wire wr_en,
	input wire clk_50m,
	input wire clken,
	output reg tx,
	output wire tx_rdy
 );

initial begin 
	tx = 1'b1;		/* Always transmit high */
end

parameter STATE_IDLE  = 2'b00;
parameter STATE_START = 2'b01;
parameter STATE_DATA  = 2'b10;
parameter STATE_STOP  = 2'b11;

reg [8:0] data = 8'h00;					// Extra parity bit
reg [3:0] bitpos = 3'h0;
reg [1:0] state = STATE_IDLE;

always @(posedge clk_50m) 
begin
	case (state)
	STATE_IDLE:
		begin
			if(wr_en)
			begin
				state <= STATE_START;	/* If write is enabled move to next state. */
				data <= din;
				bitpos <= 3'h0;
			end
		
		end
	
	STATE_START: 
	begin
			if (clken)
			begin
					tx <= 1'b0;
		   		state <= STATE_DATA;		/* Signal start by driving output to low */
			end
	end
		
	STATE_DATA:
		begin
			if (clken) 
				begin
					if (bitpos == 4'h8)
						state <= STATE_STOP;
					else
						bitpos <= bitpos + 3'h1;
					
					tx <= data[bitpos];
					
					if (bitpos < 8)
						data[8] <= data[8] ^ data[bitpos];
				end
		end
		
	STATE_STOP:
		begin
			if (clken)
				begin
					tx <= 1'b1;
					state <= STATE_IDLE;
				end
		end
		
	default:
		begin
			tx <= 1'b1;
			state <= STATE_IDLE;
		end
		
	endcase

end

assign tx_rdy = (state == STATE_IDLE);

endmodule
